library verilog;
use verilog.vl_types.all;
entity encoder8to3_vlg_vec_tst is
end encoder8to3_vlg_vec_tst;
