library verilog;
use verilog.vl_types.all;
entity demux1to4_vlg_vec_tst is
end demux1to4_vlg_vec_tst;
